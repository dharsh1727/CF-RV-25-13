
/*
See LICENSE for details
This file has been generated by CSR-BOX - 1.7.0
Time of Generation: 2025-07-24 16:37:19.466339
*/
////////////////CSR DECODER////////////////
package csrbox_decoder;
   
import Vector           :: *;
import FIFOF            :: * ;
import DReg             :: * ;
import UniqueWrappers   :: * ;
import ConcatReg        :: * ;
import GetPut           :: * ;
import Connectable      :: * ;
import csr_types        :: * ;
import Assert           :: * ;
`include "csrbox.defines"
`include "Logger.bsv"

    function Bool address_valid(Bit#(12) addr, Bit#(26) misa, Bit#(1) fs);
    Bool valid=False;
    case(addr)
   
                  `MISA:  valid= True;
                  `TDATA1: valid = True;
          	  `TDATA2: valid = True;
		  `MCONTROL6: valid = True;
                  `MVENDORID:  valid= True;
                  `STVEC: if (misa[18] == 1) valid= True;
                  `MTVEC:  valid= True;
                  `MSTATUS:  valid= True;
                  `SSTATUS: if (misa[18] == 1) valid= True;
                  `MARCHID:  valid= True;
                  `MIMPID:  valid= True;
                  `MHARTID:  valid= True;
                  `MIP:  valid= True;
                  `SIP: if (misa[18] == 1) valid= True;
                  `MIE:  valid= True;
                  `SIE: if (misa[18] == 1) valid= True;
                  `MSCRATCH:  valid= True;
                  `SSCRATCH: if (misa[18] == 1) valid= True;
                  `SEPC: if (misa[18] == 1) valid= True;
                  `STVAL: if (misa[18] == 1) valid= True;
                  `SCAUSE: if (misa[18] == 1) valid= True;
                  `MEPC:  valid= True;
                  `MTVAL:  valid= True;
                  `MCAUSE:  valid= True;
                  `MCYCLE:  valid= True;
                  `MINSTRET:  valid= True;
                  `FCSR: if (fs!=0) valid= True;
                  `TIME:  valid= True;
                  `MIDELEG:  valid= True;
                  `MEDELEG:  valid= True;
                  `PMPCFG0:  valid= True;
                  `PMPCFG2:  valid= True;
                  `PMPADDR0:  valid= True;
                  `PMPADDR1:  valid= True;
                  `PMPADDR2:  valid= True;
                  `PMPADDR3:  valid= True;
                  `PMPADDR4:  valid= True;
                  `PMPADDR5:  valid= True;
                  `PMPADDR6:  valid= True;
                  `PMPADDR7:  valid= True;
                  `PMPADDR8:  valid= True;
                  `PMPADDR9:  valid= True;
                  `PMPADDR10:  valid= True;
                  `PMPADDR11:  valid= True;
                  `PMPADDR12:  valid= True;
                  `PMPADDR13:  valid= True;
                  `PMPADDR14:  valid= True;
                  `PMPADDR15:  valid= True;
                  `MCOUNTEREN:  valid= True;
                  `SCOUNTEREN: if (misa[18] == 1) valid= True;
                  `MHPMCOUNTER3:  valid= True;
                  `MHPMCOUNTER4:  valid= True;
                  `MHPMCOUNTER5:  valid= True;
                  `MHPMCOUNTER6:  valid= True;
                  `HPMCOUNTER3:  valid= True;
                  `HPMCOUNTER4:  valid= True;
                  `HPMCOUNTER5:  valid= True;
                  `HPMCOUNTER6:  valid= True;
                  `MHPMEVENT3:  valid= True;
                  `MHPMEVENT4:  valid= True;
                  `MHPMEVENT5:  valid= True;
                  `MHPMEVENT6:  valid= True;
                  `SATP: if (misa[18] == 1) valid= True;
                  `MCOUNTINHIBIT:  valid= True;
                  `MHPMEVENT7:  valid= True;
                  `MHPMCOUNTER7:  valid= True;
                  `MHPMEVENT8:  valid= True;
                  `MHPMCOUNTER8:  valid= True;
                  `MHPMEVENT9:  valid= True;
                  `MHPMCOUNTER9:  valid= True;
                  `MHPMEVENT10:  valid= True;
                  `MHPMCOUNTER10:  valid= True;
                  `MHPMEVENT11:  valid= True;
                  `MHPMCOUNTER11:  valid= True;
                  `MHPMEVENT12:  valid= True;
                  `MHPMCOUNTER12:  valid= True;
                  `MHPMEVENT13:  valid= True;
                  `MHPMCOUNTER13:  valid= True;
                  `MHPMEVENT14:  valid= True;
                  `MHPMCOUNTER14:  valid= True;
                  `MHPMEVENT15:  valid= True;
                  `MHPMCOUNTER15:  valid= True;
                  `MHPMEVENT16:  valid= True;
                  `MHPMCOUNTER16:  valid= True;
                  `MHPMEVENT17:  valid= True;
                  `MHPMCOUNTER17:  valid= True;
                  `MHPMEVENT18:  valid= True;
                  `MHPMCOUNTER18:  valid= True;
                  `MHPMEVENT19:  valid= True;
                  `MHPMCOUNTER19:  valid= True;
                  `MHPMEVENT20:  valid= True;
                  `MHPMCOUNTER20:  valid= True;
                  `MHPMEVENT21:  valid= True;
                  `MHPMCOUNTER21:  valid= True;
                  `MHPMEVENT22:  valid= True;
                  `MHPMCOUNTER22:  valid= True;
                  `MHPMEVENT23:  valid= True;
                  `MHPMCOUNTER23:  valid= True;
                  `MHPMEVENT24:  valid= True;
                  `MHPMCOUNTER24:  valid= True;
                  `MHPMEVENT25:  valid= True;
                  `MHPMCOUNTER25:  valid= True;
                  `MHPMEVENT26:  valid= True;
                  `MHPMCOUNTER26:  valid= True;
                  `MHPMEVENT27:  valid= True;
                  `MHPMCOUNTER27:  valid= True;
                  `MHPMEVENT28:  valid= True;
                  `MHPMCOUNTER28:  valid= True;
                  `MHPMEVENT29:  valid= True;
                  `MHPMCOUNTER29:  valid= True;
                  `MHPMEVENT30:  valid= True;
                  `MHPMCOUNTER30:  valid= True;
                  `MHPMEVENT31:  valid= True;
                  `MHPMCOUNTER31:  valid= True;
                  `FFLAGS: if (fs!=0) valid= True;
                  `FRM: if (fs!=0) valid= True;
                  `CYCLE:  valid= True;
                  `INSTRET:  valid= True;
                  `HPMCOUNTER7:  valid= True;
                  `HPMCOUNTER8:  valid= True;
                  `HPMCOUNTER9:  valid= True;
                  `HPMCOUNTER10:  valid= True;
                  `HPMCOUNTER11:  valid= True;
                  `HPMCOUNTER12:  valid= True;
                  `HPMCOUNTER13:  valid= True;
                  `HPMCOUNTER14:  valid= True;
                  `HPMCOUNTER15:  valid= True;
                  `HPMCOUNTER16:  valid= True;
                  `HPMCOUNTER17:  valid= True;
                  `HPMCOUNTER18:  valid= True;
                  `HPMCOUNTER19:  valid= True;
                  `HPMCOUNTER20:  valid= True;
                  `HPMCOUNTER21:  valid= True;
                  `HPMCOUNTER22:  valid= True;
                  `HPMCOUNTER23:  valid= True;
                  `HPMCOUNTER24:  valid= True;
                  `HPMCOUNTER25:  valid= True;
                  `HPMCOUNTER26:  valid= True;
                  `HPMCOUNTER27:  valid= True;
                  `HPMCOUNTER28:  valid= True;
                  `HPMCOUNTER29:  valid= True;
                  `HPMCOUNTER30:  valid= True;
                  `HPMCOUNTER31:  valid= True;
                  `CUSTOMCONTROL:  valid= True;
                  `DCSR:  valid= True;
                  `DPC:  valid= True;
                  `DSCRATCH0:  valid= True;
                  `DSCRATCH1:  valid= True;
           endcase
     return valid;
     endfunction
    function String fn_csr_to_str(Bit#(12) addr);
    case(addr)
    
                  `MISA: return "c769_misa";
                  `MVENDORID: return "c3857_mvendorid";
                  `STVEC: return "c261_stvec";
                  `MTVEC: return "c773_mtvec";
                  `MSTATUS: return "c768_mstatus";
                  `SSTATUS: return "c256_sstatus";
                  `MARCHID: return "c3858_marchid";
                  `MIMPID: return "c3859_mimpid";
                  `MHARTID: return "c3860_mhartid";
                  `MIP: return "c836_mip";
                  `SIP: return "c324_sip";
                  `MIE: return "c772_mie";
                  `SIE: return "c260_sie";
                  `MSCRATCH: return "c832_mscratch";
                  `SSCRATCH: return "c320_sscratch";
                  `SEPC: return "c321_sepc";
                  `STVAL: return "c323_stval";
                  `SCAUSE: return "c322_scause";
                  `MEPC: return "c833_mepc";
                  `MTVAL: return "c835_mtval";
                  `MCAUSE: return "c834_mcause";
                  `MCYCLE: return "c2816_mcycle";
                  `MINSTRET: return "c2818_minstret";
                  `FCSR: return "c3_fcsr";
                  `TIME: return "c3073_time";
                  `MIDELEG: return "c771_mideleg";
                  `MEDELEG: return "c770_medeleg";
                  `PMPCFG0: return "c928_pmpcfg0";
                  `PMPCFG2: return "c930_pmpcfg2";
                  `PMPADDR0: return "c944_pmpaddr0";
                  `PMPADDR1: return "c945_pmpaddr1";
                  `PMPADDR2: return "c946_pmpaddr2";
                  `PMPADDR3: return "c947_pmpaddr3";
                  `PMPADDR4: return "c948_pmpaddr4";
                  `PMPADDR5: return "c949_pmpaddr5";
                  `PMPADDR6: return "c950_pmpaddr6";
                  `PMPADDR7: return "c951_pmpaddr7";
                  `PMPADDR8: return "c952_pmpaddr8";
                  `PMPADDR9: return "c953_pmpaddr9";
                  `PMPADDR10: return "c954_pmpaddr10";
                  `PMPADDR11: return "c955_pmpaddr11";
                  `PMPADDR12: return "c956_pmpaddr12";
                  `PMPADDR13: return "c957_pmpaddr13";
                  `PMPADDR14: return "c958_pmpaddr14";
                  `PMPADDR15: return "c959_pmpaddr15";
                  `MCOUNTEREN: return "c774_mcounteren";
                  `SCOUNTEREN: return "c262_scounteren";
                  `MHPMCOUNTER3: return "c2819_mhpmcounter3";
                  `MHPMCOUNTER4: return "c2820_mhpmcounter4";
                  `MHPMCOUNTER5: return "c2821_mhpmcounter5";
                  `MHPMCOUNTER6: return "c2822_mhpmcounter6";
                  `HPMCOUNTER3: return "c3075_hpmcounter3";
                  `HPMCOUNTER4: return "c3076_hpmcounter4";
                  `HPMCOUNTER5: return "c3077_hpmcounter5";
                  `HPMCOUNTER6: return "c3078_hpmcounter6";
                  `MHPMEVENT3: return "c803_mhpmevent3";
                  `MHPMEVENT4: return "c804_mhpmevent4";
                  `MHPMEVENT5: return "c805_mhpmevent5";
                  `MHPMEVENT6: return "c806_mhpmevent6";
                  `SATP: return "c384_satp";
                  `MCOUNTINHIBIT: return "c800_mcountinhibit";
                  `MHPMEVENT7: return "c807_mhpmevent7";
                  `MHPMCOUNTER7: return "c2823_mhpmcounter7";
                  `MHPMEVENT8: return "c808_mhpmevent8";
                  `MHPMCOUNTER8: return "c2824_mhpmcounter8";
                  `MHPMEVENT9: return "c809_mhpmevent9";
                  `MHPMCOUNTER9: return "c2825_mhpmcounter9";
                  `MHPMEVENT10: return "c810_mhpmevent10";
                  `MHPMCOUNTER10: return "c2826_mhpmcounter10";
                  `MHPMEVENT11: return "c811_mhpmevent11";
                  `MHPMCOUNTER11: return "c2827_mhpmcounter11";
                  `MHPMEVENT12: return "c812_mhpmevent12";
                  `MHPMCOUNTER12: return "c2828_mhpmcounter12";
                  `MHPMEVENT13: return "c813_mhpmevent13";
                  `MHPMCOUNTER13: return "c2829_mhpmcounter13";
                  `MHPMEVENT14: return "c814_mhpmevent14";
                  `MHPMCOUNTER14: return "c2830_mhpmcounter14";
                  `MHPMEVENT15: return "c815_mhpmevent15";
                  `MHPMCOUNTER15: return "c2831_mhpmcounter15";
                  `MHPMEVENT16: return "c816_mhpmevent16";
                  `MHPMCOUNTER16: return "c2832_mhpmcounter16";
                  `MHPMEVENT17: return "c817_mhpmevent17";
                  `MHPMCOUNTER17: return "c2833_mhpmcounter17";
                  `MHPMEVENT18: return "c818_mhpmevent18";
                  `MHPMCOUNTER18: return "c2834_mhpmcounter18";
                  `MHPMEVENT19: return "c819_mhpmevent19";
                  `MHPMCOUNTER19: return "c2835_mhpmcounter19";
                  `MHPMEVENT20: return "c820_mhpmevent20";
                  `MHPMCOUNTER20: return "c2836_mhpmcounter20";
                  `MHPMEVENT21: return "c821_mhpmevent21";
                  `MHPMCOUNTER21: return "c2837_mhpmcounter21";
                  `MHPMEVENT22: return "c822_mhpmevent22";
                  `MHPMCOUNTER22: return "c2838_mhpmcounter22";
                  `MHPMEVENT23: return "c823_mhpmevent23";
                  `MHPMCOUNTER23: return "c2839_mhpmcounter23";
                  `MHPMEVENT24: return "c824_mhpmevent24";
                  `MHPMCOUNTER24: return "c2840_mhpmcounter24";
                  `MHPMEVENT25: return "c825_mhpmevent25";
                  `MHPMCOUNTER25: return "c2841_mhpmcounter25";
                  `MHPMEVENT26: return "c826_mhpmevent26";
                  `MHPMCOUNTER26: return "c2842_mhpmcounter26";
                  `MHPMEVENT27: return "c827_mhpmevent27";
                  `MHPMCOUNTER27: return "c2843_mhpmcounter27";
                  `MHPMEVENT28: return "c828_mhpmevent28";
                  `MHPMCOUNTER28: return "c2844_mhpmcounter28";
                  `MHPMEVENT29: return "c829_mhpmevent29";
                  `MHPMCOUNTER29: return "c2845_mhpmcounter29";
                  `MHPMEVENT30: return "c830_mhpmevent30";
                  `MHPMCOUNTER30: return "c2846_mhpmcounter30";
                  `MHPMEVENT31: return "c831_mhpmevent31";
                  `MHPMCOUNTER31: return "c2847_mhpmcounter31";
                  `FFLAGS: return "c1_fflags";
                  `FRM: return "c2_frm";
                  `CYCLE: return "c3072_cycle";
                  `INSTRET: return "c3074_instret";
                  `HPMCOUNTER7: return "c3079_hpmcounter7";
                  `HPMCOUNTER8: return "c3080_hpmcounter8";
                  `HPMCOUNTER9: return "c3081_hpmcounter9";
                  `HPMCOUNTER10: return "c3082_hpmcounter10";
                  `HPMCOUNTER11: return "c3083_hpmcounter11";
                  `HPMCOUNTER12: return "c3084_hpmcounter12";
                  `HPMCOUNTER13: return "c3085_hpmcounter13";
                  `HPMCOUNTER14: return "c3086_hpmcounter14";
                  `HPMCOUNTER15: return "c3087_hpmcounter15";
                  `HPMCOUNTER16: return "c3088_hpmcounter16";
                  `HPMCOUNTER17: return "c3089_hpmcounter17";
                  `HPMCOUNTER18: return "c3090_hpmcounter18";
                  `HPMCOUNTER19: return "c3091_hpmcounter19";
                  `HPMCOUNTER20: return "c3092_hpmcounter20";
                  `HPMCOUNTER21: return "c3093_hpmcounter21";
                  `HPMCOUNTER22: return "c3094_hpmcounter22";
                  `HPMCOUNTER23: return "c3095_hpmcounter23";
                  `HPMCOUNTER24: return "c3096_hpmcounter24";
                  `HPMCOUNTER25: return "c3097_hpmcounter25";
                  `HPMCOUNTER26: return "c3098_hpmcounter26";
                  `HPMCOUNTER27: return "c3099_hpmcounter27";
                  `HPMCOUNTER28: return "c3100_hpmcounter28";
                  `HPMCOUNTER29: return "c3101_hpmcounter29";
                  `HPMCOUNTER30: return "c3102_hpmcounter30";
                  `HPMCOUNTER31: return "c3103_hpmcounter31";
                  `CUSTOMCONTROL: return "c2048_customcontrol";
                  `DCSR: return "c1968_dcsr";
                  `DPC: return "c1969_dpc";
                  `DSCRATCH0: return "c1970_dscratch0";
                  `DSCRATCH1: return "c1971_dscratch1";
                  `TDATA1: return "c1972_tdata1";
		  `TDATA2: return "c1973_tdata2";
                  `MCONTROL6: return "c1974_mcontrol6";
           endcase
     endfunction

    function Bool fn_csrbox_access(Bit#(12) csr_addr, Bit#(5) operand, Bit#(2) operation, Bit#(2) prv);
      Bool write = (operand != 0 || operation=='b01) ? True:False;
      return ((prv >= csr_addr[9:8]) && !(write && csr_addr[11:10]==2'b11) );
    endfunction:fn_csrbox_access


    
    /*doc:func: This function controls if the pipeline should be flushed for
    current csr op being decoded/processed. The control bits are used for
    dynamic control and have the following behavior: 
      - 00 : this is the default behavior where a flush is skipped for : read ops on all csrs that do not have read-side-effects (known at design time), writes on all read-only csrs
      - 01 : in this configuration a flush is skipped for only writes to on read-only csrs
      - 10 : in this configuration a flush is skipped for read-ops on all csrs do not have read-side-effects (known at design time)
      - 11 : a flush is generated for all csr ops.
    */
    function Bool fn_csr_flush(Bit#(12) addr, Bit#(3) op, Bit#(5) rs1, Bit#(2) control);

      Bool read_op = (op[1:0] == 2 || op[1:0] == 3) && rs1 == 0;
      if (control == 'b11) // flush for all read and write ops
        return True;
      else if (control[1] == 1 && !read_op ) // flush on all write ops
        return True;
      else if (control[0] == 1 && read_op) // flush on all read ops
        return True;
      else if (read_op) // do not flush on reads of any csrs
        return False;
      else // do not flush on writes to read-only csrs. Flush for all other writes
        case(addr)
        `MVENDORID , `MARCHID , `MIMPID , `MHARTID , `PMPADDR4 , `PMPADDR5 , `PMPADDR6 , `PMPADDR7 , `PMPADDR8 , `PMPADDR9 , `PMPADDR10 , `PMPADDR11 , `PMPADDR12 , `PMPADDR13 , `PMPADDR14 , `PMPADDR15 , `MCOUNTINHIBIT , `MHPMEVENT7 , `MHPMCOUNTER7 , `MHPMEVENT8 , `MHPMCOUNTER8 , `MHPMEVENT9 , `MHPMCOUNTER9 , `MHPMEVENT10 , `MHPMCOUNTER10 , `MHPMEVENT11 , `MHPMCOUNTER11 , `MHPMEVENT12 , `MHPMCOUNTER12 , `MHPMEVENT13 , `MHPMCOUNTER13 , `MHPMEVENT14 , `MHPMCOUNTER14 , `MHPMEVENT15 , `MHPMCOUNTER15 , `MHPMEVENT16 , `MHPMCOUNTER16 , `MHPMEVENT17 , `MHPMCOUNTER17 , `MHPMEVENT18 , `MHPMCOUNTER18 , `MHPMEVENT19 , `MHPMCOUNTER19 , `MHPMEVENT20 , `MHPMCOUNTER20 , `MHPMEVENT21 , `MHPMCOUNTER21 , `MHPMEVENT22 , `MHPMCOUNTER22 , `MHPMEVENT23 , `MHPMCOUNTER23 , `MHPMEVENT24 , `MHPMCOUNTER24 , `MHPMEVENT25 , `MHPMCOUNTER25 , `MHPMEVENT26 , `MHPMCOUNTER26 , `MHPMEVENT27 , `MHPMCOUNTER27 , `MHPMEVENT28 , `MHPMCOUNTER28 , `MHPMEVENT29 , `MHPMCOUNTER29 , `MHPMEVENT30 , `MHPMCOUNTER30 , `MHPMEVENT31 , `MHPMCOUNTER31 , `TDATA1, `TDATA2, `MCONTROL6 : return False;
        default: return True;
        endcase
    endfunction:fn_csr_flush


endpackage 
