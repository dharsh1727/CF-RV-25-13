
/*
See LICENSE for details
This file has been generated by CSR-BOX - 1.7.0
Time of Generation: 2025-07-24 16:37:19.498030
*/

package csrbox;
   
import Vector           :: *;
import FIFOF            :: * ;
import DReg             :: * ;
import UniqueWrappers   :: * ;
import ConcatReg        :: * ;
import GetPut           :: * ;
import Connectable      :: * ;
import csr_types        :: * ;
import Assert           :: * ;
`include "csrbox.defines"
`include "Logger.bsv"
import ccore_types :: * ;
import csrbox_grp1 :: * ;
import csrbox_grp2 :: * ;
import csrbox_decoder :: * ;
  interface Sbread;
    method Bit#(64) mv_csr_misa;
    method Bit#(32) mv_csr_mvendorid;
    method Bit#(64) mv_csr_stvec;
    method Bit#(64) mv_csr_mtvec;
    method Bit#(64) mv_csr_mstatus;
    method Bit#(64) mv_csr_marchid;
    method Bit#(64) mv_csr_mimpid;
    method Bit#(64) mv_csr_mhartid;
    method Bit#(64) mv_csr_mip;
    method Bit#(64) mv_csr_sip;
    method Bit#(64) mv_csr_mie;
    method Bit#(64) mv_csr_sie;
    method Bit#(64) mv_csr_mscratch;
    method Bit#(64) mv_csr_sscratch;
    method Bit#(64) mv_csr_sepc;
    method Bit#(64) mv_csr_stval;
    method Bit#(64) mv_csr_scause;
    method Bit#(64) mv_csr_mepc;
    method Bit#(64) mv_csr_mtval;
    method Bit#(64) mv_csr_mcause;
    method Bit#(64) mv_csr_mcycle;
    method Bit#(64) mv_csr_minstret;
    method Bit#(64) mv_csr_fcsr;
    method Bit#(64) mv_csr_time;
    method Bit#(64) mv_csr_mideleg;
    method Bit#(64) mv_csr_medeleg;
    method Bit#(64) mv_csr_pmpcfg0;
    method Bit#(30) mv_csr_pmpaddr0;
    method Bit#(30) mv_csr_pmpaddr1;
    method Bit#(30) mv_csr_pmpaddr2;
    method Bit#(30) mv_csr_pmpaddr3;
    method Bit#(32) mv_csr_mcounteren;
    method Bit#(32) mv_csr_scounteren;
    method Bit#(64) mv_csr_satp;
    method Bit#(32) mv_csr_mcountinhibit;
    method Bit#(5) mv_csr_fflags;
    method Bit#(3) mv_csr_frm;
    method Bit#(64) mv_csr_customcontrol;
    method Bit#(64) mv_csr_mhpmcounter3;
    method Bit#(64) mv_csr_mhpmcounter4;
    method Bit#(64) mv_csr_mhpmcounter5;
    method Bit#(64) mv_csr_mhpmcounter6;
    method Bit#(64) mv_csr_mhpmevent3;
    method Bit#(64) mv_csr_mhpmevent4;
    method Bit#(64) mv_csr_mhpmevent5;
    method Bit#(64) mv_csr_mhpmevent6;
    method Bit#(64) mv_csr_dcsr;
    method Bit#(64) mv_csr_dpc;
    method Bit#(64) mv_csr_dscratch0;
    method Bit#(64) mv_csr_dscratch1;

    method Bit#(64) mv_csr_tdata1;	// inserted
    method Bit#(64) mv_csr_tdata2;
    method Bit#(64) mv_csr_mcontrol6;   // inserted

  endinterface:Sbread
  // Interaface declaration
  interface Ifc_csrbox;
    interface Sbread sbread;
    method Action ma_stop_count(Bit#(1) _stop);
    method Action ma_events(Bit#(`mhpm_eventcount) events);

    method Vector#(4, Bit#(8)) mv_pmpcfg;
    method Vector#(4, Bit#(32)) mv_pmpaddr;
    method Action ma_set_mip_meip (Bit#(1) _meip);
    method Action ma_set_mip_mtip (Bit#(1) _mtip);
    method Action ma_set_mip_msip (Bit#(1) _msip);
    method Action ma_set_mip_seip (Bit#(1) _seip);
    method Action ma_incr_minstret(Bit#(64) incr);
    method Action ma_set_time (Bit#(64) _time);
    method Action ma_set_fflags (Bit#(5) _fflags, RFType rdtype);
    method Action ma_set_mip_debug_interrupt (Bit#(1) _debug_interrupt);
    method Bit#(1) mv_debug_mode;
    method Bit#(1) mv_stop_count;
    method Bit#(1) mv_stop_timer;

    
    /*doc:method : to receive the request from the core or previous node" */
    method Action ma_core_req(CSRReq req); 

    /*doc:method : to send response to core on a hit in this node" */
    method CSRResponse mv_core_resp;

    method ActionValue#(Bit#(64)) mav_upd_on_ret (Bit#(8) retype);
    
    method ActionValue#(Bit#(64)) mav_upd_on_trap(Bit#(`causesize) cause, Bit#(64) pc, Bit#(64) tval);

    method Privilege_mode mv_prv;
    
    method Bit#(1) mv_virtual;



  endinterface

  //Module Declarations
`ifdef csrbox_noinline
  (*synthesize*)
  
  (*conflict_free="ma_core_req,mv_core_resp"*)
(*conflict_free="ma_incr_minstret,sbread.mv_csr_minstret"*)
(*mutually_exclusive="mav_upd_on_trap,x0_mkConnectionAVtoAf"*)
(*mutually_exclusive="mav_upd_on_ret,x0_mkConnectionAVtoAf"*)
(*preempts="x0_mkConnectionAVtoAf,grp2_rl_increment_mhpmc3"*)
(*preempts="x0_mkConnectionAVtoAf,grp2_rl_increment_mhpmc4"*)
(*preempts="x0_mkConnectionAVtoAf,grp2_rl_increment_mhpmc5"*)
(*preempts="x0_mkConnectionAVtoAf,grp2_rl_increment_mhpmc6"*)
`endif
  module mk_csrbox(Ifc_csrbox);

    String csrbox = "";

    let grp1 <- mk_csrbox_grp1;
    let grp2 <- mk_csrbox_grp2;

    let lv_misa_s = grp1.mv_csr_misa[18];
    let lv_misa_h = grp1.mv_csr_misa[7];
    let lv_misa_u = grp1.mv_csr_misa[20];
    let lv_misa_n = grp1.mv_csr_misa[13];
    let lv_misa_c = grp1.mv_csr_misa[2];
    /*doc:reg: holds the current privilege level*/
    Reg#(Privilege_mode) rg_prv <- mkReg(Machine);
    /*doc:reg: holds the current virtual mode */
    Reg#(Bit#(1)) rg_virtual <- mkReg(0);

    /*doc:reg:The register indicates that the core is in debug mode*/
    Reg#(Bit#(1)) rg_debug_mode <- mkReg(0);

    Bool anyhit = grp1.mv_core_resp.hit || grp2.mv_core_resp.hit;
    Bit#(64) anydata = grp1.mv_core_resp.data | grp2.mv_core_resp.data;
`ifdef rtldump
    Bool anyupdated = grp1.mv_core_resp.csr_updated || grp2.mv_core_resp.csr_updated ;
`endif
    Wire#(Bit#(1)) wr_stop_count <- mkDWire(0);
    mkConnection(grp1.ma_stop_count, wr_stop_count);
    Wire#(Bit#(`mhpm_eventcount)) wr_events <- mkWire();
    mkConnection(grp2.ma_events, wr_events);
    mkConnection(grp2.ma_stop_count, wr_stop_count);

    let x0 <- mkConnection(grp1.mav_fwd_req,grp2.ma_core_req);
    mkConnection(grp1.ma_upd_privilege, rg_prv);
    mkConnection(grp1.ma_upd_virtual, rg_virtual);
    mkConnection(grp1.ma_upd_debug_mode, rg_debug_mode);
    mkConnection(grp2.ma_upd_privilege, rg_prv);
    mkConnection(grp2.ma_upd_virtual, rg_virtual);
    mkConnection(grp2.ma_upd_debug_mode, rg_debug_mode);
    mkConnection(grp2.ma_read_mcountinhibit, grp1.mv_csr_mcountinhibit);
    method mv_core_resp = CSRResponse{hit:anyhit, data: anydata 
        `ifdef rtldump , csr_updated: anyupdated `endif };
    method mv_prv = rg_prv;
    method mv_virtual = rg_virtual; 
    method ActionValue#(Bit#(64)) mav_upd_on_ret (Bit#(8) retype);
      Privilege_mode prv = unpack(retype[5:4]);
      Bool dret = (retype[3:0] == 'hb);
      Bit#(TSub#(64,1)) lv_epc = ?;

      
      if (dret) begin
        dynamicAssert(rg_debug_mode==1,"Executing DRET when not in Debug Mode");
        lv_epc = truncateLSB(grp2.mv_csr_dpc);
        rg_debug_mode <= 0;
        rg_prv <= unpack(grp2.mv_csr_dcsr[1:0]);
        if (grp2.mv_csr_dcsr[1:0] < 3)
          grp1.ma_set_mstatus_mprv(0);

      end
      else

      begin
        if (prv == Supervisor) begin
          grp1.ma_set_mstatus_spie(1'b1);
          grp1.ma_set_mstatus_sie(grp1.mv_csr_mstatus[5]);
          rg_prv <= unpack(zeroExtend(grp1.mv_csr_mstatus[8]));
          lv_epc = truncateLSB(grp1.mv_csr_sepc);
          if (lv_misa_u == 1)
            grp1.ma_set_mstatus_spp(0);
          else
            grp1.ma_set_mstatus_spp(1);
          grp1.ma_set_mstatus_mprv(0);
        end
        if (prv == Machine) begin
          rg_prv <= unpack(grp1.mv_csr_mstatus[12:11]);
          grp1.ma_set_mstatus_mpie(1'b1);
          grp1.ma_set_mstatus_mie(grp1.mv_csr_mstatus[7]);
          lv_epc = truncateLSB(grp1.mv_csr_mepc);

          if (lv_misa_u == 1)
            grp1.ma_set_mstatus_mpp(pack(User));
          else
            grp1.ma_set_mstatus_mpp(pack(Machine));

          if (grp1.mv_csr_mstatus[12:11] != '1)
            grp1.ma_set_mstatus_mprv(0);

        end
      end
      if (lv_misa_c == 0)
        lv_epc[0] = 0;
      return {lv_epc, 1'b0};
    endmethod

    method ActionValue#(Bit#(64)) mav_upd_on_trap(Bit#(`causesize) cause, Bit#(64) pc, Bit#(64) tval);
      Bit#(TSub#(`causesize,1)) lv_cause = truncate(cause);
      Bit#(1) lv_trap_type = truncateLSB(cause);
      Bit#(64) lv_tvec = ?;
      Bit#(2) lv_trapmode = 0;
      Privilege_mode prv = Machine;
      let medeleg = grp1.mv_csr_medeleg;
      let mideleg = grp1.mv_csr_mideleg;
      Bool delegateM = (truncate(mideleg >> lv_cause) & lv_trap_type) == 1 ||
                       (truncate(medeleg >> lv_cause) & ~lv_trap_type) == 1 ;
      if (delegateM && (pack(rg_prv) <= pack(Supervisor)) && lv_misa_s == 1)
        prv = Supervisor;
      
      `logLevel( csrbox, 0, $format("Taking Trap. Cause:%h,PC:%h,TVAL:%h",cause, pc, tval))
      `logLevel( csrbox, 0, $format("Trap delegated to ",fshow(prv)))

      
      if ( (lv_trap_type == 0 && (lv_cause == `halt_ebreak || 
                                lv_cause == `halt_trigger ||
                                lv_cause == `halt_step ||
                                lv_cause == `halt_reset ))
            || (lv_trap_type == 1 && lv_cause == `debug_interrupt)) begin
        grp2.ma_set_dpc(pc);
        grp2.ma_set_dcsr_cause(lv_trap_type == 1? 3:truncate(lv_cause));
        rg_debug_mode <= 1;
        grp2.ma_set_dcsr_prv(pack(rg_prv));
        rg_prv <= Machine;
        lv_tvec = `debug_parking_loop;
      end
      else if(rg_debug_mode == 1)
        lv_tvec = (lv_cause == 3 && lv_trap_type == 0)?`debug_parking_loop: `debug_parking_loop + 8;
      else

      begin

        if (prv == Supervisor) begin
          rg_prv <= Supervisor;
          grp1.ma_set_stval(tval);
          grp1.ma_set_sepc(pc);
          grp1.ma_set_scause({lv_trap_type, 'd0, lv_cause});
          grp1.ma_set_mstatus_sie(0);
          grp1.ma_set_mstatus_spp(truncate(pack(rg_prv)));
          grp1.ma_set_mstatus_spie(grp1.mv_csr_mstatus[1]);
          lv_trapmode = truncate(grp1.mv_csr_stvec);
          lv_tvec = {truncateLSB(grp1.mv_csr_stvec), 2'b0};
        end

        if (prv == Machine) begin
          rg_prv <= Machine;
          grp1.ma_set_mtval(tval);
          grp1.ma_set_mepc(pc);
          grp1.ma_set_mcause({lv_trap_type, 'd0, lv_cause});
          grp1.ma_set_mstatus_mie(1'b0);
          grp1.ma_set_mstatus_mpp(pack(rg_prv));
          grp1.ma_set_mstatus_mpie(grp1.mv_csr_mstatus[3]);
          lv_trapmode = truncate(grp1.mv_csr_mtvec);
          lv_tvec = {truncateLSB(grp1.mv_csr_mtvec), 2'b0};
        end

        if ( lv_trapmode == 1 && lv_trap_type == 1)
          lv_tvec =  lv_tvec + {zeroExtend(lv_cause),2'b0};
      end 
      `logLevel( csrbox, 0, $format("TVEC:%h",lv_tvec))
      return lv_tvec;
    endmethod
        
    method Action ma_stop_count(Bit#(1) _stop);
      wr_stop_count <= _stop;
    endmethod
    method Action ma_events(Bit#(`mhpm_eventcount) events);
      wr_events <= events;
    endmethod

    method Vector#(4, Bit#(32)) mv_pmpaddr;
        Vector#(4, Bit#(32)) lv_pmpaddr;
        lv_pmpaddr[0] = {truncate(grp1.mv_csr_pmpaddr0),2'b0};
        lv_pmpaddr[1] = {truncate(grp1.mv_csr_pmpaddr1),2'b0};
        lv_pmpaddr[2] = {truncate(grp1.mv_csr_pmpaddr2),2'b0};
        lv_pmpaddr[3] = {truncate(grp1.mv_csr_pmpaddr3),2'b0};

        return lv_pmpaddr;
    endmethod:mv_pmpaddr

    method Vector#(4, Bit#(8)) mv_pmpcfg;
        Vector#(4, Bit#(8)) lv_pmpcfg;
        lv_pmpcfg[0] = grp1.mv_csr_pmpcfg0[7:0];
        lv_pmpcfg[1] = grp1.mv_csr_pmpcfg0[15:8];
        lv_pmpcfg[2] = grp1.mv_csr_pmpcfg0[23:16];
        lv_pmpcfg[3] = grp1.mv_csr_pmpcfg0[31:24];

        return lv_pmpcfg;
    endmethod:mv_pmpcfg

    method Action ma_core_req(CSRReq req) ;
        grp1.ma_core_req(req);
    endmethod 
    interface Sbread sbread;
      method mv_csr_misa = grp1.mv_csr_misa;

      method mv_csr_mvendorid = grp1.mv_csr_mvendorid;

      method mv_csr_stvec = grp1.mv_csr_stvec;

      method mv_csr_mtvec = grp1.mv_csr_mtvec;

      method mv_csr_mstatus = grp1.mv_csr_mstatus;

      method mv_csr_marchid = grp1.mv_csr_marchid;

      method mv_csr_mimpid = grp1.mv_csr_mimpid;

      method mv_csr_mhartid = grp1.mv_csr_mhartid;

      method mv_csr_mip = grp1.mv_csr_mip;

      method mv_csr_sip = grp1.mv_csr_sip;

      method mv_csr_mie = grp1.mv_csr_mie;

      method mv_csr_sie = grp1.mv_csr_sie;

      method mv_csr_mscratch = grp1.mv_csr_mscratch;

      method mv_csr_sscratch = grp1.mv_csr_sscratch;

      method mv_csr_sepc = grp1.mv_csr_sepc;

      method mv_csr_stval = grp1.mv_csr_stval;

      method mv_csr_scause = grp1.mv_csr_scause;

      method mv_csr_mepc = grp1.mv_csr_mepc;

      method mv_csr_mtval = grp1.mv_csr_mtval;

      method mv_csr_mcause = grp1.mv_csr_mcause;

      method mv_csr_mcycle = grp1.mv_csr_mcycle;

      method mv_csr_minstret = grp1.mv_csr_minstret;

      method mv_csr_fcsr = grp1.mv_csr_fcsr;

      method mv_csr_time = grp1.mv_csr_time;

      method mv_csr_mideleg = grp1.mv_csr_mideleg;

      method mv_csr_medeleg = grp1.mv_csr_medeleg;

      method mv_csr_pmpcfg0 = grp1.mv_csr_pmpcfg0;

      method mv_csr_pmpaddr0 = grp1.mv_csr_pmpaddr0;

      method mv_csr_pmpaddr1 = grp1.mv_csr_pmpaddr1;

      method mv_csr_pmpaddr2 = grp1.mv_csr_pmpaddr2;

      method mv_csr_pmpaddr3 = grp1.mv_csr_pmpaddr3;

      method mv_csr_mcounteren = grp1.mv_csr_mcounteren;

      method mv_csr_scounteren = grp1.mv_csr_scounteren;

      method mv_csr_satp = grp1.mv_csr_satp;

      method mv_csr_mcountinhibit = grp1.mv_csr_mcountinhibit;

      method mv_csr_fflags = grp1.mv_csr_fflags;

      method mv_csr_frm = grp1.mv_csr_frm;

      method mv_csr_customcontrol = grp1.mv_csr_customcontrol;

      method mv_csr_mhpmcounter3 = grp2.mv_csr_mhpmcounter3;

      method mv_csr_mhpmcounter4 = grp2.mv_csr_mhpmcounter4;

      method mv_csr_mhpmcounter5 = grp2.mv_csr_mhpmcounter5;

      method mv_csr_mhpmcounter6 = grp2.mv_csr_mhpmcounter6;

      method mv_csr_mhpmevent3 = grp2.mv_csr_mhpmevent3;

      method mv_csr_mhpmevent4 = grp2.mv_csr_mhpmevent4;

      method mv_csr_mhpmevent5 = grp2.mv_csr_mhpmevent5;

      method mv_csr_mhpmevent6 = grp2.mv_csr_mhpmevent6;

      method mv_csr_dcsr = grp2.mv_csr_dcsr;

      method mv_csr_dpc = grp2.mv_csr_dpc;

      method mv_csr_dscratch0 = grp2.mv_csr_dscratch0;

      method mv_csr_dscratch1 = grp2.mv_csr_dscratch1;
      
      method mv_csr_tdata1 = grp2.mv_csr_tdata1;	 //inserted
      method mv_csr_tdata2 = grp2.mv_csr_tdata2;
      method mv_csr_mcontrol6 = grp2.mv_csr_mcontrol6;   //inserted

    endinterface
    method ma_set_mip_meip = grp1.ma_set_mip_meip;
    method ma_set_mip_mtip = grp1.ma_set_mip_mtip;
    method ma_set_mip_msip = grp1.ma_set_mip_msip;
    method ma_set_mip_seip = grp1.ma_set_mip_seip;
    method ma_incr_minstret = grp1.ma_incr_minstret;
    method ma_set_time = grp1.ma_set_time;
    method ma_set_fflags = grp1.ma_set_fflags;
    method ma_set_mip_debug_interrupt = grp1.ma_set_mip_debug_interrupt;
    method mv_debug_mode = rg_debug_mode;
    method mv_stop_count = pack(rg_debug_mode) & grp2.mv_csr_dcsr[10];
    method mv_stop_timer = pack(rg_debug_mode) & grp2.mv_csr_dcsr[9];

  endmodule 
endpackage 
