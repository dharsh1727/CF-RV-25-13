
/*
See LICENSE for details
This file has been generated by CSR-BOX - 1.7.0
Time of Generation: 2025-07-28 21:04:28.315704
*/

package csr_types ;
    `include "csrbox.defines"
    `include "Logger.bsv"


    typedef struct {
        Bit#(12) csr_address;
        Bit#(64) writedata;
        Bit#(2) funct3;
        Bit#(1) pc_1;
    } CSRReq deriving(Bits, FShow, Eq);

    typedef struct{
        Bool hit;
        Bit#(64)  data;
    `ifdef rtldump
        Bool csr_updated;
    `endif
    } CSRResponse deriving(Bits, Eq, FShow);
    
    // -----------------------------------------------
    // Trigger-related types for mcontrol6-style trigger
    // -----------------------------------------------

    typedef struct {
        Bit#(32) tdata1;
        Bit#(32) tdata2;
    } TriggerData0 deriving (Bits, FShow);
    
  typedef struct {
    Bit#(4)   type_t;        // bits [3:0]
    Bit#(1)   dmode;       // bit [4]
    Bit#(6)   maskmax;     // bits [10:5]
    Bit#(2)   sizehi;      // bits [12:11]
    Bit#(1)   select;      // bit [13]
    Bit#(1)   timing;      // bit [14]
    Bit#(2)   size;        // bits [16:15]
    Bit#(4)   action_;      // bits [20:17]
    Bit#(1)   chain;       // bit [21]
    Bit#(4)   match_type;  // bits [25:22]
    Bit#(1)   machine;     // bit [26]
    Bit#(1)   supervisor;  // bit [27]
    Bit#(1)   user;        // bit [28]
    Bit#(1)   execute;     // bit [29]
    Bit#(1)   store;       // bit [30]
    Bit#(1)   load;        // bit [31]
  } Mcontrol6 deriving (Bits, Eq, FShow);
    typedef enum {Machine = 3, Hypervisor=2, Supervisor = 1, User = 0} Privilege_mode deriving(Bits, Eq, FShow);


    function Bit#(64) fn_csr_op (Bit#(64) writedata, Bit#(64) readdata, Bit#(2) op);
        if(op == 'd1)
    	    return writedata;
        else if(op == 'd2)
            return (writedata|readdata);
        else
            return (~writedata & readdata);
    endfunction
  
  function Reg#(Bit#(1)) extInterruptReg(Reg#(Bit#(1)) r1, Reg#(Bit#(1)) r2);
    return (interface Reg;
      method Bit#(1) _read = r1 | r2;
      method Action _write(Bit#(1) x);
        r1._write(x);
      endmethod
    endinterface);
  endfunction
  
endpackage 
