
/*
See LICENSE for details
This file has been generated by CSR-BOX - 1.7.0
Time of Generation: 2025-07-28 21:04:28.344813
*/

package csrbox_grp2;
   
import Vector           :: *;
import FIFOF            :: * ;
import DReg             :: * ;
import UniqueWrappers   :: * ;
import ConcatReg        :: * ;
import GetPut           :: * ;
import Connectable      :: * ;
import csr_types        :: * ;
import Assert           :: * ;
`include "csrbox.defines"
`include "Logger.bsv"
import ccore_types :: * ;

  // Interaface declaration
  interface Ifc_csrbox_grp2;
    method Action ma_events(Bit#(`mhpm_eventcount) events);
    method Action ma_stop_count(Bit#(1) _stop);

    method Bit#(64) mv_csr_mhpmcounter3;
    method Bit#(64) mv_csr_mhpmcounter4;
    method Bit#(64) mv_csr_mhpmcounter5;
    method Bit#(64) mv_csr_mhpmcounter6;
    method Bit#(64) mv_csr_mhpmevent3;
    method Bit#(64) mv_csr_mhpmevent4;
    method Bit#(64) mv_csr_mhpmevent5;
    method Bit#(64) mv_csr_mhpmevent6;
    method Bit#(64) mv_csr_dcsr;
    method Bit#(64) mv_csr_dpc;
    method Bit#(64) mv_csr_dscratch0;
    method Bit#(64) mv_csr_dscratch1;

    method Bit#(64) mv_csr_tdata1;                 /*inserted*/
    method Bit#(64) mv_csr_tdata2;                 /*inserted*/
    method Mcontrol6 mv_csr_mcontrol6;             /*inserted*/   
    method TriggerData0 mv_trigger_data; 
    method Action mav_upd_on_trigger(Bit#(7) cause, Bit#(64) pc);

    
    method Action ma_set_dcsr_cause (Bit#(3) _cause);
    method Action ma_set_dcsr_prv (Bit#(2) _prv);
    method Action ma_set_dpc (Bit#(64) _dpc);


    method Action ma_read_mcountinhibit (Bit#(32) _mcountinhibit);    
    /*doc:method : to receive the request from the core or previous node" */
    method Action ma_core_req(CSRReq req); 

    /*doc:method : to send response to core on a hit in this node" */
    method CSRResponse mv_core_resp;

    /*doc:method: fetch from core the prvilege mode */
    method Action ma_upd_privilege (Privilege_mode prv);
    
    /*doc:method: fetch from core the virtual mode */
    method Action ma_upd_virtual (Bit#(1) _virtual);
    
    method Action ma_upd_debug_mode (Bit#(1) _dbg);
    
  endinterface

  //Module Declarations
`ifdef csrbox_grp_noinline
  (*synthesize*)
  
  (*conflict_free="ma_core_req,mv_core_resp"*)
  (*preempts = "ma_core_req, rl_increment_mhpmc3"*)
  (*preempts = "ma_core_req, rl_increment_mhpmc4"*)
  (*preempts = "ma_core_req, rl_increment_mhpmc5"*)
  (*preempts = "ma_core_req, rl_increment_mhpmc6"*)
  (*mutually_exclusive = "ma_set_dcsr_prv, ma_core_req"*)
  (*mutually_exclusive = "ma_set_dcsr_cause, ma_core_req"*)
  (*mutually_exclusive = "ma_set_dpc, ma_core_req"*)

`endif
  module mk_csrbox_grp2(Ifc_csrbox_grp2);

    String csrbox = "";
    Wire#(Bit#(64)) wr_mtvec <- mkWire(); 

    /*doc:wire: holds the response of this group for a csr operation request,
    for one cycle, wire is used for low latency*/
    Wire#(CSRResponse) rg_resp_to_core <- mkDWire(CSRResponse{hit:False, data:0
        `ifdef rtldump , csr_updated: False `endif });

    /*doc:fifo: fifo to forward the core request to the next group on a miss*/
    FIFOF#(CSRReq) ff_fwd_request <- mkFIFOF();

    /*doc:wire: holds the current privilege mode of the hart*/
    Wire#(Privilege_mode) wr_prv <- mkWire();
   
    /*doc:wire: holds the current state of the vs bit of the hart*/
    Wire#(Bit#(1)) wr_virtual <- mkWire();

    Wire#(Bit#(1)) wr_debug_mode <- mkWire();

    Wire#(Bit#(`mhpm_eventcount)) wr_events <- mkWire();
    Wire#(Bit#(1)) wr_stop_count <- mkDWire(0);
    /*doc:wire: */
    Wire#(Bit#(32)) rg_mcountinhibit <- mkDWire(0);

    function Reg#(Bit#(64)) warlReg_mhpmcounter3(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mhpmcounter3

    /*doc:reg: The mhpmcounter3 is a 64-bit counter. Returns lower 32 bits in RV32I mode.*/
    Reg#(Bit#(64)) rg_mhpmcounter3_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_mhpmcounter3 = warlReg_mhpmcounter3(rg_mhpmcounter3_warl);
    
    function Reg#(Bit#(64)) warlReg_tdata1(Reg#(Bit#(64)) r);			/*inserted*/
           return (interface Reg;				
                method Bit#(64) _read = r;
                method Action _write(Bit#(64) x);
                  Mcontrol6 val = unpack(truncate(x));
                  val.type_t = 6;
                  val.dmode = 1;
                  r._write(zeroExtend(pack(val)));
               endmethod
           endinterface);
    endfunction: warlReg_tdata1
 
    Reg#(Bit#(64)) rg_tdata1_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_tdata1 = warlReg_tdata1(rg_tdata1_warl);                  /*inserted*/

    function Reg#(Bit#(64)) warlReg_tdata2(Reg#(Bit#(64)) r);			/*inserted*/
            return (interface Reg;
                 method Bit#(64) _read = r;
                 method Action _write(Bit#(64) x);
                      r._write(x);
                 endmethod
            endinterface);
    endfunction: warlReg_tdata2

    Reg#(Bit#(64)) rg_tdata2_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_tdata2 = warlReg_tdata2(rg_tdata2_warl);			//inserted
    
    function Reg#(Bit#(64)) warlReg_mhpmcounter4(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mhpmcounter4

    /*doc:reg: The mhpmcounter4 is a 64-bit counter. Returns lower 42 bits in RV42I mode.*/
    Reg#(Bit#(64)) rg_mhpmcounter4_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_mhpmcounter4 = warlReg_mhpmcounter4(rg_mhpmcounter4_warl);

    function Reg#(Bit#(64)) warlReg_mhpmcounter5(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mhpmcounter5

    /*doc:reg: The mhpmcounter5 is a 64-bit counter. Returns lower 52 bits in RV52I mode.*/
    Reg#(Bit#(64)) rg_mhpmcounter5_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_mhpmcounter5 = warlReg_mhpmcounter5(rg_mhpmcounter5_warl);

    function Reg#(Bit#(64)) warlReg_mhpmcounter6(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mhpmcounter6

    /*doc:reg: The mhpmcounter6 is a 64-bit counter. Returns lower 62 bits in RV62I mode.*/
    Reg#(Bit#(64)) rg_mhpmcounter6_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_mhpmcounter6 = warlReg_mhpmcounter6(rg_mhpmcounter6_warl);

    function Reg#(Bit#(64)) warlReg_mhpmevent3(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (( x[63:0] >= 0 && x[63:0] <= 31 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mhpmevent3

    /*doc:reg: The mhpmevent3 is a MXLEN-bit event register which controls mhpmcounter3.*/
    Reg#(Bit#(64)) rg_mhpmevent3_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_mhpmevent3 = warlReg_mhpmevent3(rg_mhpmevent3_warl);

    function Reg#(Bit#(64)) warlReg_mhpmevent4(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (( x[63:0] >= 0 && x[63:0] <= 31 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mhpmevent4

    /*doc:reg: The mhpmevent4 is a MXLEN-bit event register which controls mhpmcounter4.*/
    Reg#(Bit#(64)) rg_mhpmevent4_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_mhpmevent4 = warlReg_mhpmevent4(rg_mhpmevent4_warl);

    function Reg#(Bit#(64)) warlReg_mhpmevent5(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (( x[63:0] >= 0 && x[63:0] <= 31 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mhpmevent5

    /*doc:reg: The mhpmevent5 is a MXLEN-bit event register which controls mhpmcounter5.*/
    Reg#(Bit#(64)) rg_mhpmevent5_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_mhpmevent5 = warlReg_mhpmevent5(rg_mhpmevent5_warl);

    function Reg#(Bit#(64)) warlReg_mhpmevent6(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (( x[63:0] >= 0 && x[63:0] <= 31 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_mhpmevent6

    /*doc:reg: The mhpmevent6 is a MXLEN-bit event register which controls mhpmcounter6.*/
    Reg#(Bit#(64)) rg_mhpmevent6_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_mhpmevent6 = warlReg_mhpmevent6(rg_mhpmevent6_warl);

    function Reg#(Bit#(2)) warlReg_dcsr_prv(Reg#(Bit#(2)) r);
        return (interface Reg;
            method Bit#(2) _read = r;
            method Action _write(Bit#(2) x);
               if (True) begin
                   if (( x[1:0] == 0 || x[1:0] == 1 || x[1:0] == 3 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_dcsr_prv

    /*doc:reg: Contains the privilege level the hart was operating in when Debug Mode was entered.*/
    Reg#(Bit#(2)) rg_dcsr_prv_warl <- mkReg(3);
    Reg#(Bit#(2)) rg_dcsr_prv = warlReg_dcsr_prv(rg_dcsr_prv_warl);

    function Reg#(Bit#(1)) warlReg_dcsr_step(Reg#(Bit#(1)) r);
        return (interface Reg;
            method Bit#(1) _read = r;
            method Action _write(Bit#(1) x);
               if (True) begin
                   if (( x[0] == 0 || x[0] == 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_dcsr_step

    /*doc:reg: When set and not in Debug Mode the hart will only execute a single instruction;then enter Debug Mode*/
    Reg#(Bit#(1)) rg_dcsr_step_warl <- mkReg(0);
    Reg#(Bit#(1)) rg_dcsr_step = warlReg_dcsr_step(rg_dcsr_step_warl);

    /*doc:reg: When set, there is a Non-Maskable-Interrupt (NMI) pending for the hart.*/
    Reg#(Bit#(1)) rg_dcsr_nmip <- mkReg(0);

    function Reg#(Bit#(1)) warlReg_dcsr_mprven(Reg#(Bit#(1)) r);
        return (interface Reg;
            method Bit#(1) _read = r;
            method Action _write(Bit#(1) x);
               if (True) begin
                   if (( x[0] == 0 || x[0] == 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_dcsr_mprven

    /*doc:reg: mprv in mstatus.*/
    Reg#(Bit#(1)) rg_dcsr_mprven_warl <- mkReg(0);
    Reg#(Bit#(1)) rg_dcsr_mprven = warlReg_dcsr_mprven(rg_dcsr_mprven_warl);

    /*doc:reg: Extends the prv field with the virtualization mode WARL 0 the hart was operating in when Debug Mode was entered*/
    Reg#(Bit#(1)) rg_dcsr_v = readOnlyReg(0);

    /*doc:reg: Explains why Debug Mode was entered*/
    Reg#(Bit#(3)) rg_dcsr_cause <- mkReg(0);

    function Reg#(Bit#(1)) warlReg_dcsr_stoptime(Reg#(Bit#(1)) r);
        return (interface Reg;
            method Bit#(1) _read = r;
            method Action _write(Bit#(1) x);
               if (True) begin
                   if (( x[0] == 0 || x[0] == 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_dcsr_stoptime

    /*doc:reg: Don’t increment any hart-local timers while in Debug Mode.*/
    Reg#(Bit#(1)) rg_dcsr_stoptime_warl <- mkReg(0);
    Reg#(Bit#(1)) rg_dcsr_stoptime = warlReg_dcsr_stoptime(rg_dcsr_stoptime_warl);

    function Reg#(Bit#(1)) warlReg_dcsr_stopcount(Reg#(Bit#(1)) r);
        return (interface Reg;
            method Bit#(1) _read = r;
            method Action _write(Bit#(1) x);
               if (True) begin
                   if (( x[0] == 0 || x[0] == 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_dcsr_stopcount

    /*doc:reg: Don’t increment any hart-local counters while in Debug Mode*/
    Reg#(Bit#(1)) rg_dcsr_stopcount_warl <- mkReg(0);
    Reg#(Bit#(1)) rg_dcsr_stopcount = warlReg_dcsr_stopcount(rg_dcsr_stopcount_warl);

    function Reg#(Bit#(1)) warlReg_dcsr_stepie(Reg#(Bit#(1)) r);
        return (interface Reg;
            method Bit#(1) _read = r;
            method Action _write(Bit#(1) x);
               if (True) begin
                   if (( x[0] == 0 || x[0] == 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_dcsr_stepie

    /*doc:reg: Interrupts (including NMI) are enabled during single stepping.*/
    Reg#(Bit#(1)) rg_dcsr_stepie_warl <- mkReg(0);
    Reg#(Bit#(1)) rg_dcsr_stepie = warlReg_dcsr_stepie(rg_dcsr_stepie_warl);

    function Reg#(Bit#(1)) warlReg_dcsr_ebreaku(Reg#(Bit#(1)) r);
        return (interface Reg;
            method Bit#(1) _read = r;
            method Action _write(Bit#(1) x);
               if (True) begin
                   if (( x[0] == 0 || x[0] == 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_dcsr_ebreaku

    /*doc:reg: ebreak instructions in U-mode enter Debug Mode.*/
    Reg#(Bit#(1)) rg_dcsr_ebreaku_warl <- mkReg(0);
    Reg#(Bit#(1)) rg_dcsr_ebreaku = warlReg_dcsr_ebreaku(rg_dcsr_ebreaku_warl);

    function Reg#(Bit#(1)) warlReg_dcsr_ebreaks(Reg#(Bit#(1)) r);
        return (interface Reg;
            method Bit#(1) _read = r;
            method Action _write(Bit#(1) x);
               if (True) begin
                   if (( x[0] == 0 || x[0] == 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_dcsr_ebreaks

    /*doc:reg: ebreak instructions in S-mode enter Debug Mode.*/
    Reg#(Bit#(1)) rg_dcsr_ebreaks_warl <- mkReg(0);
    Reg#(Bit#(1)) rg_dcsr_ebreaks = warlReg_dcsr_ebreaks(rg_dcsr_ebreaks_warl);

    function Reg#(Bit#(1)) warlReg_dcsr_ebreakm(Reg#(Bit#(1)) r);
        return (interface Reg;
            method Bit#(1) _read = r;
            method Action _write(Bit#(1) x);
               if (True) begin
                   if (( x[0] == 0 || x[0] == 1 )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_dcsr_ebreakm

    /*doc:reg: ebreak instructions in M-mode enter Debug Mode.*/
    Reg#(Bit#(1)) rg_dcsr_ebreakm_warl <- mkReg(0);
    Reg#(Bit#(1)) rg_dcsr_ebreakm = warlReg_dcsr_ebreakm(rg_dcsr_ebreakm_warl);

    /*doc:reg: ebreak instructions in VU-mode enter Debug Mode.*/
    Reg#(Bit#(1)) rg_dcsr_ebreakvu = readOnlyReg(0);

    /*doc:reg: ebreak instructions in VS-mode enter Debug Mode.*/
    Reg#(Bit#(1)) rg_dcsr_ebreakvs = readOnlyReg(0);

    /*doc:reg: Debug support exists as it is described in this document.*/
    Reg#(Bit#(4)) rg_dcsr_debugver = readOnlyReg(4);

    /*doc:reg: The mstatus register keeps track of and controls the hart’s current operating state. */
    Reg#(Bit#(64)) rg_dcsr = concatReg18(  readOnlyReg(32'd0) ,rg_dcsr_debugver , readOnlyReg(10'd0) ,rg_dcsr_ebreakvs ,rg_dcsr_ebreakvu ,rg_dcsr_ebreakm , readOnlyReg(1'd0) ,rg_dcsr_ebreaks ,rg_dcsr_ebreaku ,rg_dcsr_stepie ,rg_dcsr_stopcount ,rg_dcsr_stoptime ,readOnlyReg(rg_dcsr_cause), rg_dcsr_v ,rg_dcsr_mprven ,readOnlyReg(rg_dcsr_nmip), rg_dcsr_step ,rg_dcsr_prv );

    function Reg#(Bit#(64)) warlReg_dpc(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_dpc

    /*doc:reg: Upon entry to debug mode, dpc is updated with the virtual address of the next instruction to be executed.*/
    Reg#(Bit#(64)) rg_dpc_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_dpc = warlReg_dpc(rg_dpc_warl);

    function Reg#(Bit#(64)) warlReg_dscratch0(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_dscratch0

    /*doc:reg: The dscratch0 register is an DXLEN-bit read/write register dedicated for use by debug mode.*/
    Reg#(Bit#(64)) rg_dscratch0_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_dscratch0 = warlReg_dscratch0(rg_dscratch0_warl);

    function Reg#(Bit#(64)) warlReg_dscratch1(Reg#(Bit#(64)) r);
        return (interface Reg;
            method Bit#(64) _read = r;
            method Action _write(Bit#(64) x);
               if (True) begin
                   if (( True )) begin
                       let _x = x;
        
                       r._write(_x);
                   end
               end

            endmethod
        endinterface);
    endfunction: warlReg_dscratch1

    /*doc:reg: The dscratch1 register is an DXLEN-bit read/write register dedicated for use by debug mode.*/
    Reg#(Bit#(64)) rg_dscratch1_warl <- mkReg(0);
    Reg#(Bit#(64)) rg_dscratch1 = warlReg_dscratch1(rg_dscratch1_warl);
    rule rl_increment_mhpmc3;
      if (wr_stop_count == 0)
        rg_mhpmcounter3 <= rg_mhpmcounter3 + zeroExtend(~rg_mcountinhibit[3]&wr_events[rg_mhpmevent3]);
    endrule
    rule rl_increment_mhpmc4;
      if (wr_stop_count == 0)
      rg_mhpmcounter4 <= rg_mhpmcounter4 + zeroExtend(~rg_mcountinhibit[4]&wr_events[rg_mhpmevent4]);
    endrule
    rule rl_increment_mhpmc5;
      if (wr_stop_count == 0)
      rg_mhpmcounter5 <= rg_mhpmcounter5 + zeroExtend(~rg_mcountinhibit[5]&wr_events[rg_mhpmevent5]);
    endrule
    rule rl_increment_mhpmc6;
      if (wr_stop_count == 0)
      rg_mhpmcounter6 <= rg_mhpmcounter6 + zeroExtend(~rg_mcountinhibit[6]&wr_events[rg_mhpmevent6]);
    endrule
 
    method Action ma_core_req(CSRReq req);
        `logLevel( csrbox_grp2, 1, $format("csrbox_grp2: received req: ", fshow(req)))
        Bit#(2) op = req.funct3; 
        case (req.csr_address) 
            `MHPMCOUNTER3 : begin
                Bit#(64) readdata = zeroExtend(rg_mhpmcounter3);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mhpmcounter3 <= truncate(word);
            end
	    
	    `TDATA1 : begin					 /*inserted*/
                Bit#(64) readdata = rg_tdata1;
                rg_resp_to_core <= CSRResponse { hit: True, data: readdata
                           `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, req.funct3);
		rg_tdata1 <= truncate(word);
	    end							 /*inserted*/

	    `TDATA2 : begin					 /*inserted*/
  		Bit#(64) readdata = zeroExtend(rg_tdata2);
  		rg_resp_to_core <= CSRResponse { hit: True, data: readdata
    			`ifdef rtldump ,csr_updated: True `endif };
  		let word = fn_csr_op(req.writedata, readdata, req.funct3);
  		
  		rg_tdata2 <= truncate(word);

            end							 /*inserted*/
            
            `MCONTROL6: begin                                    /*inserted*/
 		 Bit#(64) readdata = zeroExtend(rg_tdata1);
  		 rg_resp_to_core <= CSRResponse { hit: True,data: readdata
    			`ifdef rtldump ,csr_updated: False `endif };
		 let word = fn_csr_op(req.writedata, readdata, req.funct3);
  		 rg_tdata1 <= truncate(word);

	     end
	     
            `MHPMCOUNTER4 : begin
                Bit#(64) readdata = zeroExtend(rg_mhpmcounter4);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mhpmcounter4 <= truncate(word);
            end

            `MHPMCOUNTER5 : begin
                Bit#(64) readdata = zeroExtend(rg_mhpmcounter5);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mhpmcounter5 <= truncate(word);
            end

            `MHPMCOUNTER6 : begin
                Bit#(64) readdata = zeroExtend(rg_mhpmcounter6);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mhpmcounter6 <= truncate(word);
            end
            `HPMCOUNTER3 : begin
                Bit#(64) readdata = truncate(rg_mhpmcounter3);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump ,csr_updated: True `endif };
            end
            `HPMCOUNTER4 : begin
                Bit#(64) readdata = truncate(rg_mhpmcounter4);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump ,csr_updated: True `endif };
            end
            `HPMCOUNTER5 : begin
                Bit#(64) readdata = truncate(rg_mhpmcounter5);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump ,csr_updated: True `endif };
            end
            `HPMCOUNTER6 : begin
                Bit#(64) readdata = truncate(rg_mhpmcounter6);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata `ifdef rtldump ,csr_updated: True `endif };
            end

            `MHPMEVENT3 : begin
                Bit#(64) readdata = zeroExtend(rg_mhpmevent3);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mhpmevent3 <= truncate(word);
            end

            `MHPMEVENT4 : begin
                Bit#(64) readdata = zeroExtend(rg_mhpmevent4);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mhpmevent4 <= truncate(word);
            end

            `MHPMEVENT5 : begin
                Bit#(64) readdata = zeroExtend(rg_mhpmevent5);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mhpmevent5 <= truncate(word);
            end

            `MHPMEVENT6 : begin
                Bit#(64) readdata = zeroExtend(rg_mhpmevent6);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_mhpmevent6 <= truncate(word);
            end

            `DCSR : begin
                Bit#(64) readdata = zeroExtend(rg_dcsr);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_dcsr <= truncate(word);
            end

            `DPC : begin
                Bit#(64) readdata = zeroExtend(rg_dpc);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_dpc <= truncate(word);
            end

            `DSCRATCH0 : begin
                Bit#(64) readdata = zeroExtend(rg_dscratch0);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_dscratch0 <= truncate(word);
            end

            `DSCRATCH1 : begin
                Bit#(64) readdata = zeroExtend(rg_dscratch1);
                rg_resp_to_core <= CSRResponse{hit:True, data: readdata
                    `ifdef rtldump ,csr_updated: True `endif };
                let word = fn_csr_op(req.writedata, readdata, op);
                
                 rg_dscratch1 <= truncate(word);
            end

            default: begin
                rg_resp_to_core <= CSRResponse{hit: True, data: 0 `ifdef rtldump , csr_updated : False `endif };
            end
        endcase
        endmethod
     
        
    method mv_csr_mhpmcounter3 = rg_mhpmcounter3;

    method mv_csr_mhpmcounter4 = rg_mhpmcounter4;

    method mv_csr_mhpmcounter5 = rg_mhpmcounter5;

    method mv_csr_mhpmcounter6 = rg_mhpmcounter6;

    method mv_csr_mhpmevent3 = rg_mhpmevent3;

    method mv_csr_mhpmevent4 = rg_mhpmevent4;

    method mv_csr_mhpmevent5 = rg_mhpmevent5;

    method mv_csr_mhpmevent6 = rg_mhpmevent6;

    method mv_csr_dcsr = rg_dcsr;

    method mv_csr_dpc = rg_dpc;

    method mv_csr_dscratch0 = rg_dscratch0;
    
    method Bit#(64) mv_csr_tdata1 = rg_tdata1;
    method Bit#(64) mv_csr_tdata2 = rg_tdata2;
    method Mcontrol6 mv_csr_mcontrol6 = unpack(truncate(rg_tdata1));

    method TriggerData0 mv_trigger_data();
        return TriggerData0 {
            tdata1: truncate(rg_tdata1),
            tdata2: truncate(rg_tdata2)
        };
    endmethod
    
    method Action mav_upd_on_trigger(Bit#(7) cause, Bit#(64) pc);
	  rg_dpc_warl <= pc;
	  rg_dcsr_cause <= truncate(pack(cause)[2:0]);
    endmethod

    method mv_csr_dscratch1 = rg_dscratch1;
    method Action ma_set_dcsr_cause (Bit#(3) _cause);
      rg_dcsr_cause <= _cause;
    endmethod
    method Action ma_set_dcsr_prv (Bit#(2) _prv);
      rg_dcsr_prv <= _prv;
    endmethod
    method Action ma_set_dpc (Bit#(64) _dpc);
      rg_dpc <= _dpc;
    endmethod

    method Action ma_read_mcountinhibit (Bit#(32) _mcountinhibit);
        rg_mcountinhibit <= _mcountinhibit;
    endmethod
    method Action ma_events(Bit#(`mhpm_eventcount) events);
      wr_events <= events;
    endmethod
    method Action ma_stop_count(Bit#(1) _stop);
      wr_stop_count <= _stop;
    endmethod

    method mv_core_resp = rg_resp_to_core;

    method Action ma_upd_privilege (Privilege_mode prv);
        wr_prv <= prv;
    endmethod
    
    method Action ma_upd_virtual (Bit#(1) _virtual);
         wr_virtual <= _virtual;
    endmethod
    method Action ma_upd_debug_mode (Bit#(1) _dbg);
        wr_debug_mode <= _dbg;
    endmethod
  endmodule 
endpackage 
