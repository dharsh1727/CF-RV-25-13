
/*
See LICENSE for details
This file has been generated by CSR-BOX - 1.7.0
Time of Generation: 2025-07-28 21:04:28.315704
*/

package csr_types ;
    `include "csrbox.defines"
    `include "Logger.bsv"


    typedef struct {
        Bit#(12) csr_address;
        Bit#(64) writedata;
        Bit#(2) funct3;
        Bit#(1) pc_1;
    } CSRReq deriving(Bits, FShow, Eq);

    typedef struct{
        Bool hit;
        Bit#(64)  data;
    `ifdef rtldump
        Bool csr_updated;
    `endif
    } CSRResponse deriving(Bits, Eq, FShow);
    
    // -----------------------------------------------
    // Trigger-related types for mcontrol6-style trigger
    // -----------------------------------------------

    typedef struct {
        Bit#(32) tdata1;
        Bit#(32) tdata2;
    } TriggerData0 deriving (Bits, FShow);
    
  typedef struct {
    Bit#(4)   type_t;        
    Bit#(1)   dmode;       
    Bit#(6)   maskmax;     
    Bit#(2)   sizehi;      
    Bit#(1)   select;
    Bit#(1)   timing;    
    Bit#(2)   size;     
    Bit#(4)   action_;      
    Bit#(1)   chain;       
    Bit#(4)   match_type;  
    Bit#(1)   machine;     
    Bit#(1)   supervisor;  
    Bit#(1)   user;        
    Bit#(1)   execute;    
    Bit#(1)   store;       
    Bit#(1)   load;        
  } Mcontrol6 deriving (Bits, Eq, FShow);
    typedef enum {Machine = 3, Hypervisor=2, Supervisor = 1, User = 0} Privilege_mode deriving(Bits, Eq, FShow);


    function Bit#(64) fn_csr_op (Bit#(64) writedata, Bit#(64) readdata, Bit#(2) op);
        if(op == 'd1)
    	    return writedata;
        else if(op == 'd2)
            return (writedata|readdata);
        else
            return (~writedata & readdata);
    endfunction
  
  function Reg#(Bit#(1)) extInterruptReg(Reg#(Bit#(1)) r1, Reg#(Bit#(1)) r2);
    return (interface Reg;
      method Bit#(1) _read = r1 | r2;
      method Action _write(Bit#(1) x);
        r1._write(x);
      endmethod
    endinterface);
  endfunction
  
endpackage 
